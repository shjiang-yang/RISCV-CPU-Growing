//================================================
//designer: shjiang
//data: 2020-06-20
//
//description:
//to decode the part of intruction in IFU
//
//===============================================

module ifu_miniDec(
    pass
)

